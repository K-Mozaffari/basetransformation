
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use WORK.Package_Moduli_Set_4_w2.ALL;

ENTITY CPA_WITH_IEAC IS ---(2^n+1)
GENERIC(n:INTEGER:=3);
PORT (Xin,Yin:IN   STD_LOGIC_VECTOR(n-1 DOWNTO 0);Cin:IN STD_LOGIC;
      Sout   :OUT  STD_LOGIC_VECTOR(n DOWNTO 0)
      );
END CPA_WITH_IEAC;

ARCHITECTURE STRUCTURAL OF CPA_WITH_IEAC IS
SIGNAL S,Sm :STD_LOGIC_VECTOR(n-1 DOWNTO 0);
SIGNAL C,C_NOT,Cm:STD_LOGIC;
BEGIN

CPAF    :CPA_FA       GENERIC MAP(n)  PORT MAP(Xin,Yin,Cin,S,C);
C_NOT<=NOT(C);
CPAH    :CPA_HA       GENERIC MAP(n)  PORT MAP(S,C_NOT,Sm,Cm);
SOUT<=Cm&Sm; 

END STRUCTURAL;