library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.package_Constant.all;
use WORK.Package_Moduli_Set_4_w2.ALL;

ENTITY BASE_TRANSFORMATION_M4_W2 IS 
  GENERIC (n:INTEGER:=4;
           a:INTEGER:=2;
           m:INTEGER:=1;
           RQ1:INTEGER:=1;
           R2:INTEGER:=1;
           R3:INTEGER:=1;
           rQ1_4:INTEGER:=1;
           R2_4:INTEGER:=1;
           R3_4:INTEGER:=1
         );
 PORT (x1_in :IN  STD_LOGIC_VECTOR(n     DOWNTO 0);
       x2_in :IN  STD_LOGIC_VECTOR(2*n-1   DOWNTO 0);
       x3_in :IN  STD_LOGIC_VECTOR(n-1   DOWNTO 0);
       x4_in :IN  STD_LOGIC_VECTOR(2*n  DOWNTO 0);
       x1_out:OUT STD_LOGIC_VECTOR(n-a   DOWNTO 0);
       x2_out:OUT STD_LOGIC_VECTOR(2*n-a-1 DOWNTO 0);
       x3_out:OUT STD_LOGIC_VECTOR(n-a-1 DOWNTO 0);
       x4_out:OUT STD_LOGIC_VECTOR(2*(n-a) DOWNTO 0)
       );
END BASE_TRANSFORMATION_M4_W2;

ARCHITECTURE STRUCTURAL OF BASE_TRANSFORMATION_M4_W2 IS 
   SIGNAL  P1,P2,P31,P32,P_S:STD_LOGIC_VECTOR(2*n-1 DOWNTO 0);
   SIGNAL  B1_S,B2_S,B3_S,BL_S:STD_LOGIC_VECTOR(m-1 DOWNTO 0);
   SIGNAL  Cp_S,SIGN:STD_LOGIC;
   SIGNAL  Q1 :STD_LOGIC_VECTOR(2*n   DOWNTO 0);
   SIGNAL  Q2 :STD_LOGIC_VECTOR(m+(4*n)-1 DOWNTO 0);
   SIGNAL  Q3 :STD_LOGIC_VECTOR(m-1 DOWNTO 0);
   SIGNAL  Sx1,Cx1,Sx3,Cx3:STD_LOGIC_VECTOR(n-a-1 DOWNTO 0);
   SIGNAL  Sx4,Cx4:STD_LOGIC_VECTOR(2*(n-a)-1 DOWNTO 0);

  BEGIN 
  
     OPU1   :OPU_1    GENERIC MAP (n)   PORT MAP (x1_in,x3_in,x4_in,P1,P2,P31,P32);
     UNITPCP:UNIT_PCp GENERIC MAP (n)   PORT MAP (P1,P2,P31,P32,P_S,Cp_S);

     OPU2   :OPU_2    GENERIC MAP (n,m) PORT MAP (P_S,x2_in,x4_in,B1_S,B2_S,B3_S);
     UNITBL :UNIT_BL  GENERIC MAP (m)   PORT MAP (B1_S,B2_S,B3_S,Cp_S,BL_S);

     OPU3   :OPU_3     GENERIC MAP(n,m ) PORT MAP (x4_in,P_S,BL_S,Q1,Q2,Q3,SIGN);

     Gx1:CSA_IEAC_TREE       GENERIC MAP (n,a,m,RQ1,R2,R3) PORT MAP (Q1,Q2,Q3,Sx1,Cx1);
     GY1:ADDER_MAPPING_IEAC  GENERIC MAP (n,a)             PORT MAP (Sx1,Cx1,RF1_BIN,C1_SIGN,C1_CARRY,C1_SIGN_CARRY,Cp_S,SIGN,x1_out);

     Gx3:CSA_EAC_TREE      GENERIC MAP (n,a,m,RQ1,R2,R3) PORT MAP (Q1,Q2,Q3,Sx3,Cx3);
     GY3:ADDER_MAPPING_EAC GENERIC MAP (n,a)             PORT MAP (Sx3,Cx3,C3_SIGN,C3_CARRY,C3_SIGN_CARRY,Cp_S,SIGN,x3_out);

     Gx4:CSA_IEAC2_TREE       GENERIC MAP (n,a,m,rQ1_4,R2_4,R3_4) PORT MAP (Q1,Q2,Q3,Sx4,Cx4);
     GY4:ADDER_MAPPING_IEAC2  GENERIC MAP (n,a)                   PORT MAP (Sx4,Cx4,RF4_BIN,C4_SIGN,C4_CARRY,C4_SIGN_CARRY,Cp_S,SIGN,x4_out);
x2_out<=x2_in(2*n-a-1 DOWNTO 0);

END STRUCTURAL;
