

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use WORK.Package_Moduli_Set_4_w2.ALL;

ENTITY OPU_1 IS 
 GENERIC (n:INTEGER:=5 );
 PORT (x1 :IN  STD_LOGIC_VECTOR(n     DOWNTO 0);
       x3 :IN  STD_LOGIC_VECTOR(n-1   DOWNTO 0);
       x4 :IN  STD_LOGIC_VECTOR(2*n   DOWNTO 0);
       P1 :OUT STD_LOGIC_VECTOR(2*n-1 DOWNTO 0);
       P2 :OUT STD_LOGIC_VECTOR(2*n-1 DOWNTO 0);
       P31:OUT STD_LOGIC_VECTOR(2*n-1 DOWNTO 0);
       P32:OUT STD_LOGIC_VECTOR(2*n-1 DOWNTO 0)
      );
END OPU_1;

ARCHITECTURE STRUCTURAL OF OPU_1 IS
  SIGNAL x1_NOT:STD_LOGIC_VECTOR(n   DOWNTO 0);
  SIGNAL x4_NOT:STD_LOGIC_VECTOR(2*n DOWNTO 0);
  SIGNAL VDD   :STD_LOGIC_VECTOR(n-3 DOWNTO 0):=(OTHERS=>'1');
  SIGNAL GND   :STD_LOGIC_VECTOR(n-2 DOWNTO 0):=(OTHERS=>'0');
 BEGIN
   x1_NOT<=NOT(x1);
   x4_NOT<=NOT(x4);
   P1 <=x1(1)&x1(0)&GND   (n-2   DOWNTO 0)&x1 (n   DOWNTO 2);
   P2 <=x3(1)&x3(0)&x3    (n-1   DOWNTO 0)&x3 (n-1 DOWNTO 2);
   P31<=x4_NOT(2*n)&x1_NOT(n     DOWNTO 0)&VDD(n-3 DOWNTO 0);
   P32<=x4_NOT(0)  &x4_NOT(2*n-1 DOWNTO 1);
END STRUCTURAL;


