
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use WORK.Package_Moduli_Set_4_w2.ALL;

ENTITY CPA_WITH_EAC IS ---(2^2n-1)
 GENERIC(n:INTEGER:=2);
 PORT (Xin,Yin:IN   STD_LOGIC_VECTOR(n-1 DOWNTO 0);
       Sout   :OUT  STD_LOGIC_VECTOR(n-1 DOWNTO 0)
       );
END CPA_WITH_EAC;

ARCHITECTURE STRUCTURAL OF CPA_WITH_EAC IS
  SIGNAL S :STD_LOGIC_VECTOR(n-1 DOWNTO 0);
  SIGNAL C,D,DC:STD_LOGIC;
  SIGNAL GND:STD_LOGIC:='0';
 BEGIN
  CPAF    :CPA_FA       GENERIC MAP(n)  PORT MAP(Xin,Yin,GND,S,C);
  DETECTOR:DETECTOR_ONE GENERIC MAP(n)  PORT MAP(S,D);
  DC<=D OR C;
  CPAH    :CPA_HA       GENERIC MAP(n)  PORT MAP(S,DC,Sout,OPEN);
END STRUCTURAL;