
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use WORK.Package_Moduli_Set_4_w2.ALL;

ENTITY UNIT_PCp is---(Adder 2^2n-1)
 GENERIC (n : INTEGER := 3
	 );
	PORT (	P1_in : IN  STD_LOGIC_VECTOR(2*n-1 DOWNTO 0);
		P2_in : IN  STD_LOGIC_VECTOR(2*n-1 DOWNTO 0);
		P31_in: IN  STD_LOGIC_VECTOR(2*n-1 DOWNTO 0);
		P32_in: IN  STD_LOGIC_VECTOR(2*n-1 DOWNTO 0);
		P_out : OUT STD_LOGIC_VECTOR(2*n-1 DOWNTO 0);
		Cp    : OUT STD_LOGIC
	      );
END UNIT_PCp;

ARCHITECTURE STRUCTURAL OF UNIT_PCp IS 
   SIGNAL S2,C2,S1,C1,Sm:STD_LOGIC_VECTOR(2*n-1 DOWNTO 0);
   SIGNAL D             :STD_LOGIC;
   SIGNAL GND           :STD_LOGIC_VECTOR(2*n-1 DOWNTO 0):=(OTHERS=>'0');
  BEGIN
   CSA1   :CSA_WITH_EAC  GENERIC MAP (2*n) PORT MAP(P1_in,P2_in,P31_in,S1,C1);
   CSA2   :CSA_WITH_EAC  GENERIC MAP (2*n) PORT MAP(S1 ,C1 ,P32_in,S2 ,C2 );  
   CPA    :CPA_FA        GENERIC MAP (2*n) PORT MAP(S2 ,C2,GND(0) ,Sm,Cp);
   DETECTE:DETECTOR_ONE  GENERIC MAP (2*n) PORT MAP (Sm,D);
   MUX:mux2to1           GENERIC MAP (2*n) port map (Sm,GND,D,P_out);
  END STRUCTURAL;
