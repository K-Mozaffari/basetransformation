library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
package Package_Constant is
CONSTANT n:integer:=8;
CONSTANT a:integer:=2;
CONSTANT Rif:integer:=6;
CONSTANT C1:STD_LOGIC_VECTOR(n-a-1 DOWNTO 0):="111010";
CONSTANT C2:STD_LOGIC_VECTOR(n-a-1 DOWNTO 0):="111100";
CONSTANT C3:STD_LOGIC_VECTOR(2*(n-a)-1 DOWNTO 0):="000001000010";
END PACKAGE;