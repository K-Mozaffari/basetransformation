library IEEE;

use IEEE.STD_LOGIC_1164.ALL;
use work.package_Constant.all;
use work.Package_Moduli_Set_4_w2.all;

ENTITY ADDER_MAPPING_EAC IS
 GENERIC (n:INTEGER:=4;
          a:INTEGER:=2
           );   
 PORT (Sx3          :IN  STD_LOGIC_VECTOR(n-a-1 DOWNTO 0);
       Cx3          :IN  STD_LOGIC_VECTOR(n-a-1 DOWNTO 0);
       C3_SIGN      :IN  STD_LOGIC_VECTOR(n-a-1 DOWNTO 0);
       C3_CARRY     :IN  STD_LOGIC_VECTOR(n-a-1 DOWNTO 0);
       C3_SIGN_CARRY:IN  STD_LOGIC_VECTOR(n-a-1 DOWNTO 0);
       Cp           :IN  STD_LOGIC;
       SIGN         :IN  STD_LOGIC;
       x_3          :OUT STD_LOGIC_VECTOR(n-a-1 DOWNTO 0)
       );
	    
END ADDER_MAPPING_EAC;

ARCHITECTURE STRUCTURAL OF ADDER_MAPPING_EAC IS
   SIGNAL S1,C1,OMUX:STD_LOGIC_VECTOR(n-a-1 DOWNTO 0);
   SIGNAL GND:STD_LOGIC_VECTOR(n-a-1 DOWNTO 0):=(OTHERS=>'0');
   SIGNAL SEL:STD_LOGIC_VECTOR(1 DOWNTO 0);
 BEGIN 
SEL<=Cp&SIGN;
   MUX:MUX4TO1       GENERIC MAP (n-a) PORT MAP (GND,C3_SIGN,C3_CARRY,C3_SIGN_CARRY,SEL,OMUX);   
   CSA:CSA_WITH_EAC  GENERIC MAP (n-a) PORT MAP (Sx3,Cx3,OMUX,S1,C1); 
   CPA:CPA_WITH_EAC  GENERIC MAP (n-a) PORT MAP (S1,C1,x_3);
END STRUCTURAL;

