
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use WORK.Package_Moduli_Set_4_w2.ALL;

ENTITY UNIT_BL is---(Adder 2^n)
 GENERIC (n : INTEGER := 3
	  );
 PORT    (	B1_in : IN  STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		B2_in : IN  STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		B3_in : IN  STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		Cp    : IN  STD_LOGIC;
		BL_out: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0)
	  );
END UNIT_BL;

ARCHITECTURE STRUCTURAL OF UNIT_BL IS 
   SIGNAL S1,C1,S2,C2,Dc   :std_logic_vector(n-1 DOWNTO 0);
   SIGNAL VDD:STD_LOGIC:='1';
   SIGNAL GND:STD_LOGIC_VECTOR(n-2 DOWNTO 0):=(OTHERS=>'0');
  BEGIN
Dc<=GND(n-2 DOWNTO 0)&Cp;
   CSA_1  :CSA    GENERIC MAP(n)    PORT MAP(B1_in,B2_in,B3_in,S1,C1);
   CSA_2  :CSA    GENERIC MAP(n)    PORT MAP(S1,C1,Dc,S2,C2);
   CPA    :CPA_FA             GENERIC MAP(n)    PORT MAP(S2,C2,VDD,BL_out,OPEN);
END STRUCTURAL;
